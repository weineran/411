/* cache.sv
 *	The cache design. It contains the cache controller and cache datapath.
 */
 